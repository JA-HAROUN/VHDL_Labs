LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY test_Ripple IS
END test_Ripple;

ARCHITECTURE tbRippleAdder OF test_Ripple IS

    COMPONENT RippleAdder IS
        PORT (
            A_3 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            B_3 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            CarryIn : IN STD_LOGIC;
            Sum : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            CarryOut : OUT STD_LOGIC
        );
    END COMPONENT;

    SIGNAL A, B : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
    SIGNAL Cin : STD_LOGIC := '0';
    SIGNAL S : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL Cout : STD_LOGIC;

BEGIN

    R : RippleAdder PORT MAP(
        A_3 => A,
        B_3 => B,
        CarryIn => Cin,
        Sum => S,
        CarryOut => Cout
    );

    PROCESS BEGIN

        WAIT FOR 2 ns;

        FOR i IN 0 TO 1 LOOP

            FOR j IN 0 TO 15 LOOP

                FOR k IN 0 TO 15 LOOP

                    -- change A
                    A <= STD_LOGIC_VECTOR(unsigned(A) + 1);
                    WAIT FOR 1 ns;

                END LOOP;

                -- change B
                B <= STD_LOGIC_VECTOR(unsigned(B) + 1);
                WAIT FOR 1 ns;

            END LOOP;

            -- change Cin
            Cin <= NOT Cin;
            WAIT FOR 1 ns;

        END LOOP;

        WAIT;

    END PROCESS;

END tbRippleAdder;